case 16h0000: { mem_rdata = 0xC001; }
case 16h0001: { mem_rdata = 0xC000; }
case 16h0002: { mem_rdata = 0x97FF; }
case 16h0003: { mem_rdata = 0x9531; }
case 16h0004: { mem_rdata = 0xA522; }
case 16h0005: { mem_rdata = 0x9811; }
case 16h0006: { mem_rdata = 0xA80A; }
case 16h0007: { mem_rdata = 0x6582; }
case 16h0008: { mem_rdata = 0x4758; }
case 16h0009: { mem_rdata = 0x82FE; }
case 16h000A: { mem_rdata = 0x6585; }
case 16h000B: { mem_rdata = 0x4758; }
case 16h000C: { mem_rdata = 0x6585; }
case 16h000D: { mem_rdata = 0x4758; }
case 16h000E: { mem_rdata = 0x6820; }
case 16h000F: { mem_rdata = 0x6520; }
case 16h0010: { mem_rdata = 0x4758; }
case 16h0011: { mem_rdata = 0xC102; }
case 16h0012: { mem_rdata = 0x0302; }
case 16h0013: { mem_rdata = 0xD003; }
case 16h0014: { mem_rdata = 0xFFFF; }
case 16h0015: { mem_rdata = 0x0007; }
