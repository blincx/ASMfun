case 16h0000: { mem_rdata = 0xC001; }
case 16h0001: { mem_rdata = 0xC000; }
case 16h0002: { mem_rdata = 0x8802; }
case 16h0003: { mem_rdata = 0x8B03; }
case 16h0004: { mem_rdata = 0x97FF; }
case 16h0005: { mem_rdata = 0x68B2; }
case 16h0006: { mem_rdata = 0x0E1D; }
case 16h0007: { mem_rdata = 0x9CFF; }
case 16h0008: { mem_rdata = 0xACFC; }
case 16h0009: { mem_rdata = 0x8502; }
case 16h000A: { mem_rdata = 0x061A; }
case 16h000B: { mem_rdata = 0x0517; }
case 16h000C: { mem_rdata = 0x8A00; }
case 16h000D: { mem_rdata = 0x8801; }
case 16h000E: { mem_rdata = 0x6680; }
case 16h000F: { mem_rdata = 0x4960; }
case 16h0010: { mem_rdata = 0xD009; }
case 16h0011: { mem_rdata = 0xFFFF; }
case 16h0012: { mem_rdata = 0x8A30; }
case 16h0013: { mem_rdata = 0x47A8; }
case 16h0014: { mem_rdata = 0xD005; }
case 16h0015: { mem_rdata = 0x8A31; }
case 16h0016: { mem_rdata = 0x47A8; }
case 16h0017: { mem_rdata = 0xD005; }
case 16h0018: { mem_rdata = 0x8A32; }
case 16h0019: { mem_rdata = 0x47A8; }
case 16h001A: { mem_rdata = 0xD005; }
case 16h001B: { mem_rdata = 0x8A33; }
case 16h001C: { mem_rdata = 0x47A8; }
case 16h001D: { mem_rdata = 0xD005; }
case 16h001E: { mem_rdata = 0x47A8; }
case 16h001F: { mem_rdata = 0x47C8; }
case 16h0020: { mem_rdata = 0x6C50; }
case 16h0021: { mem_rdata = 0xD20E; }
case 16h0022: { mem_rdata = 0xFFFF; }
case 16h0023: { mem_rdata = 0x000C; }
case 16h0024: { mem_rdata = 0x000A; }
case 16h0025: { mem_rdata = 0x0026; }
case 16h0026: { mem_rdata = 0x0012; }
case 16h0027: { mem_rdata = 0x0015; }
case 16h0028: { mem_rdata = 0x0018; }
case 16h0029: { mem_rdata = 0x001B; }
case 16h002A: { mem_rdata = 0x001E; }
